
.global gnd vdd

*** TOP LEVEL CELL: Inverter{sch}
Mnmos@1 out in gnd gnd NMOS L=0.4U W=4U
Mpmos@1 vdd in out vdd PMOS L=0.4U W=2U

* Spice Code nodes in cell cell 'Inverter{sch}'
vdd vdd 0 DC 5
vin in 0 DC pwl 10n 0 20n 5 50n 5 60n 0
cload out 0 250fF
.measure tran tf trig v(out) val=4.5 fall=1 td=8ns targ v(out) val=0.5 fall=1
.measure tran tr trig v(out) val=0.5 rise=1 td=50ns targ v(out) val=4.5 rise=1
.tran 0 100n
*.dc vin 0 5 1m
.include C:\Users\Vaasudeva\Documents\electric\180nm2.txt
.END
