
.global gnd vdd

*** TOP LEVEL CELL: sram:sram{sch}
Mnmos@0 gnd q qb gnd NMOS L=0.4U W=2U
Mnmos@1 q qb gnd gnd NMOS L=0.4U W=2U
Mnmos@2 qb wl bl gnd NMOS L=0.4U W=2U
Mnmos@3 blb wl q gnd NMOS L=0.4U W=2U
Mpmos@0 qb q vdd vdd PMOS L=0.4U W=2U
Mpmos@1 vdd qb q vdd PMOS L=0.4U W=2U

* Spice Code nodes in cell cell 'sram:sram{sch}'
vdd vdd 0 dc 5
vwl wl 0 dc pwl 10n 0 20n 5 50n 5 60n 5 90n 5 100n 0 130n 0 140n 0 170n 0 180n 5
vbl bl 0 dc pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vblb blb 0 dc pwl 10n 5 20n 0 50n 0 60n 5 90n 5 100n 0 130n 0 140n 5 170n 5 180n 0
.tran 0 200n
.include C:\Users\Vaasudeva\Documents\electric\180nm2.txt
.END
