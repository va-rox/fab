
*** TOP LEVEL CELL: sram:sram_lay{lay}
Mnmos@0 q qb net@8 gnd NMOS L=0.4U W=2U AS=43.62P AD=3.62P PS=35.4U PD=11.4U
Mnmos@1 net@8 q qb gnd NMOS L=0.4U W=2U AS=3.62P AD=43.62P PS=11.4U PD=35.4U
Mnmos@2 q wl bl gnd NMOS L=0.4U W=2U AS=9.62P AD=3.62P PS=25.4U PD=11.4U
Mnmos@3 blb wl qb gnd NMOS L=0.4U W=2U AS=3.62P AD=9.62P PS=11.4U PD=25.4U
Mpmos@0 q qb net@4 vdd PMOS L=0.4U W=2U AS=43.62P AD=3.62P PS=35.4U PD=11.4U
Mpmos@1 net@4 q qb vdd PMOS L=0.4U W=2U AS=3.62P AD=43.62P PS=11.4U PD=35.4U

* Spice Code nodes in cell cell 'sram:sram_lay{lay}'
vdd vdd 0 dc 5
vwl wl 0 dc pwl 10n 0 20n 5 50n 5 60n 5 90n 5 100n 0 130n 5 140n 0 170n 0 180n 5
vbl bl 0 dc pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vblb blb 0 dc pwl 10n 5 20n 0 50n 0 60n 5 90n 5 100n 0 130n 0 140n 5 170n 5 180n 0
.tran 0 200n
.include C:\Users\Vaasudeva\Documents\electric\180nm2.txt
.END
